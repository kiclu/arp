library verilog;
use verilog.vl_types.all;
entity shftr32_vlg_vec_tst is
end shftr32_vlg_vec_tst;
