library verilog;
use verilog.vl_types.all;
entity mx4_32b_vlg_vec_tst is
end mx4_32b_vlg_vec_tst;
