library verilog;
use verilog.vl_types.all;
entity reg32_ld_clr_vlg_vec_tst is
end reg32_ld_clr_vlg_vec_tst;
