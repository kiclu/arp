library verilog;
use verilog.vl_types.all;
entity dc3_8_vlg_vec_tst is
end dc3_8_vlg_vec_tst;
