library verilog;
use verilog.vl_types.all;
entity cmp32s_vlg_vec_tst is
end cmp32s_vlg_vec_tst;
