library verilog;
use verilog.vl_types.all;
entity rv32i_vlg_vec_tst is
end rv32i_vlg_vec_tst;
