library verilog;
use verilog.vl_types.all;
entity gpu_vlg_vec_tst is
end gpu_vlg_vec_tst;
