library verilog;
use verilog.vl_types.all;
entity shftl32_vlg_vec_tst is
end shftl32_vlg_vec_tst;
