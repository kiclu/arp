library verilog;
use verilog.vl_types.all;
entity reg1_ld_clr_vlg_vec_tst is
end reg1_ld_clr_vlg_vec_tst;
