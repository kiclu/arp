library verilog;
use verilog.vl_types.all;
entity regfile_vlg_vec_tst is
end regfile_vlg_vec_tst;
