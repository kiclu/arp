library verilog;
use verilog.vl_types.all;
entity pc_vlg_vec_tst is
end pc_vlg_vec_tst;
