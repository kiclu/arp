library verilog;
use verilog.vl_types.all;
entity dram_init_vlg_vec_tst is
end dram_init_vlg_vec_tst;
