library verilog;
use verilog.vl_types.all;
entity dc2_4_vlg_vec_tst is
end dc2_4_vlg_vec_tst;
