library verilog;
use verilog.vl_types.all;
entity mx2_32b_vlg_vec_tst is
end mx2_32b_vlg_vec_tst;
