library verilog;
use verilog.vl_types.all;
entity reg11_ld_clr_inc_vlg_vec_tst is
end reg11_ld_clr_inc_vlg_vec_tst;
