library verilog;
use verilog.vl_types.all;
entity cmp4_vlg_vec_tst is
end cmp4_vlg_vec_tst;
