library verilog;
use verilog.vl_types.all;
entity reg16_ld_clr_vlg_vec_tst is
end reg16_ld_clr_vlg_vec_tst;
