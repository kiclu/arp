library verilog;
use verilog.vl_types.all;
entity shftl_vlg_vec_tst is
end shftl_vlg_vec_tst;
