library verilog;
use verilog.vl_types.all;
entity sram_controller_vlg_vec_tst is
end sram_controller_vlg_vec_tst;
