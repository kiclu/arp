library verilog;
use verilog.vl_types.all;
entity cmp4_vlg_check_tst is
    port(
        E1              : in     vl_logic;
        G1              : in     vl_logic;
        L1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end cmp4_vlg_check_tst;
