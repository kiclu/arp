library verilog;
use verilog.vl_types.all;
entity dif_vlg_vec_tst is
end dif_vlg_vec_tst;
