library verilog;
use verilog.vl_types.all;
entity vga_hfp_vlg_check_tst is
    port(
        vga_hfp         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end vga_hfp_vlg_check_tst;
