library verilog;
use verilog.vl_types.all;
entity reg8_ld_clr_vlg_vec_tst is
end reg8_ld_clr_vlg_vec_tst;
