library verilog;
use verilog.vl_types.all;
entity reg1_ld_clr_vlg_check_tst is
    port(
        DOUT            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end reg1_ld_clr_vlg_check_tst;
