library verilog;
use verilog.vl_types.all;
entity ARP_vlg_vec_tst is
end ARP_vlg_vec_tst;
