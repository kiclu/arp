library verilog;
use verilog.vl_types.all;
entity shft16l32_vlg_vec_tst is
end shft16l32_vlg_vec_tst;
